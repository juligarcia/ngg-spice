TEMP TITLE
RR1 node-5 gnd 10K
VV1 gnd node-5 10
.tran 10u 10
.end
