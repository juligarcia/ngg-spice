TEMP TITLE
RR1 node-4 gnd 10K
VV1 node-4 gnd 10
.op
.end
