TEMP TITLE
RR1 gnd node-5 10K
VV1 gnd node-5 10
.op
.end
