TEMP TITLE
RR1 gnd node-4 10K
VV1 gnd node-4 10
.op
.end
