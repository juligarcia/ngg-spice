TEMP TITLE
RR1 node-4 gnd 10K
VV1 node-4 gnd 10
.tran 10u 10
.end
