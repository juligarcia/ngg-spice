TEMP TITLE
.tran 10u 10
.end
