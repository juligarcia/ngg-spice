TEMP TITLE
.op
.end
