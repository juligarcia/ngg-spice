TEMP TITLE
RR1 node-4 gnd 10K
VV1 gnd node-4 10
.tran 10u 10
.end
