TEMP TITLE
.end
